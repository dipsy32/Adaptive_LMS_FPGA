module rom_data (
    input wire clk,
    input wire [9:0] addr,
    output reg [31:0] data
);

    always @(posedge clk) begin
        case(addr)
            10'd0: data <= 32'h00120024;
            10'd1: data <= 32'hff9bff17;
            10'd2: data <= 32'h006fffe7;
            10'd3: data <= 32'h0030ffee;
            10'd4: data <= 32'h0080001c;
            10'd5: data <= 32'h00b2008f;
            10'd6: data <= 32'h0039ffa6;
            10'd7: data <= 32'h00b2ffd9;
            10'd8: data <= 32'h00e30075;
            10'd9: data <= 32'h0062ff92;
            10'd10: data <= 32'h01010026;
            10'd11: data <= 32'h007effa3;
            10'd12: data <= 32'h0103001d;
            10'd13: data <= 32'h0088ffa8;
            10'd14: data <= 32'h00ecfffe;
            10'd15: data <= 32'h0074ff7c;
            10'd16: data <= 32'h015b00e9;
            10'd17: data <= 32'h0076003d;
            10'd18: data <= 32'h00b1000f;
            10'd19: data <= 32'h00940029;
            10'd20: data <= 32'h003fff9f;
            10'd21: data <= 32'h0026ff48;
            10'd22: data <= 32'h00820018;
            10'd23: data <= 32'h001afff7;
            10'd24: data <= 32'hfff7ffa1;
            10'd25: data <= 32'hfff3ffb5;
            10'd26: data <= 32'h000f0033;
            10'd27: data <= 32'hff9cffc3;
            10'd28: data <= 32'hffadffbd;
            10'd29: data <= 32'hff56ff5a;
            10'd30: data <= 32'hffff008e;
            10'd31: data <= 32'hff9300b0;
            10'd32: data <= 32'hff1bffaf;
            10'd33: data <= 32'hff68ffe9;
            10'd34: data <= 32'hff0dff96;
            10'd35: data <= 32'hff20ff7d;
            10'd36: data <= 32'hff70003c;
            10'd37: data <= 32'hff5d0085;
            10'd38: data <= 32'hff390045;
            10'd39: data <= 32'hff1affdd;
            10'd40: data <= 32'hff12ff8e;
            10'd41: data <= 32'hff700016;
            10'd42: data <= 32'hff06ff86;
            10'd43: data <= 32'hff9a0017;
            10'd44: data <= 32'hff13ff6b;
            10'd45: data <= 32'hffb8fff3;
            10'd46: data <= 32'hff77ffd1;
            10'd47: data <= 32'hfff50053;
            10'd48: data <= 32'hffda005a;
            10'd49: data <= 32'h000a0067;
            10'd50: data <= 32'hfffc002d;
            10'd51: data <= 32'h0005ffe4;
            10'd52: data <= 32'hfffaff7c;
            10'd53: data <= 32'h000aff38;
            10'd54: data <= 32'h0077ffc9;
            10'd55: data <= 32'h0098003c;
            10'd56: data <= 32'h001eff46;
            10'd57: data <= 32'h00bdffc3;
            10'd58: data <= 32'h00bf002a;
            10'd59: data <= 32'h0089ffb0;
            10'd60: data <= 32'h00bbffbb;
            10'd61: data <= 32'h00ec002f;
            10'd62: data <= 32'h0079ff7b;
            10'd63: data <= 32'h00d5ffb6;
            10'd64: data <= 32'h00adffbc;
            10'd65: data <= 32'h011e008d;
            10'd66: data <= 32'h00a90041;
            10'd67: data <= 32'h00cb0041;
            10'd68: data <= 32'h0027ff3d;
            10'd69: data <= 32'h00bbffdc;
            10'd70: data <= 32'h0046ffb5;
            10'd71: data <= 32'h0051ffa3;
            10'd72: data <= 32'h008d0061;
            10'd73: data <= 32'hfff9ffce;
            10'd74: data <= 32'h0065005e;
            10'd75: data <= 32'h00130076;
            10'd76: data <= 32'hffe9002c;
            10'd77: data <= 32'hff87ff84;
            10'd78: data <= 32'hffdafffe;
            10'd79: data <= 32'hff8ffffc;
            10'd80: data <= 32'hff6cffbb;
            10'd81: data <= 32'hffb4005c;
            10'd82: data <= 32'hff660049;
            10'd83: data <= 32'hff3fffe9;
            10'd84: data <= 32'hff34ffc8;
            10'd85: data <= 32'hff81006a;
            10'd86: data <= 32'hfe75fec3;
            10'd87: data <= 32'hffb20024;
            10'd88: data <= 32'hff20003a;
            10'd89: data <= 32'hff62004c;
            10'd90: data <= 32'hff14ffe1;
            10'd91: data <= 32'hff4dffe8;
            10'd92: data <= 32'hff4ffff6;
            10'd93: data <= 32'hffb5009e;
            10'd94: data <= 32'hff28ffca;
            10'd95: data <= 32'hfff0008d;
            10'd96: data <= 32'hff56ffe1;
            10'd97: data <= 32'hffbbffd2;
            10'd98: data <= 32'hffd80012;
            10'd99: data <= 32'hffcfffdb;
            10'd100: data <= 32'hffd5ff8f;
            10'd101: data <= 32'h006d006e;
            10'd102: data <= 32'h000a0002;
            10'd103: data <= 32'h002fffa9;
            10'd104: data <= 32'h0036ff82;
            10'd105: data <= 32'h0067ff9e;
            10'd106: data <= 32'h0053ff66;
            10'd107: data <= 32'h00d20017;
            10'd108: data <= 32'h004dff68;
            10'd109: data <= 32'h012c0077;
            10'd110: data <= 32'h0081ffea;
            10'd111: data <= 32'h00defff2;
            10'd112: data <= 32'h00e00037;
            10'd113: data <= 32'h008cff9c;
            10'd114: data <= 32'h00f40011;
            10'd115: data <= 32'h00b00000;
            10'd116: data <= 32'h00cb0014;
            10'd117: data <= 32'h0094ffe3;
            10'd118: data <= 32'h010b00c3;
            10'd119: data <= 32'h00760052;
            10'd120: data <= 32'h005fffd6;
            10'd121: data <= 32'h004dffc2;
            10'd122: data <= 32'h0030ffad;
            10'd123: data <= 32'h004e000d;
            10'd124: data <= 32'hffc9ff75;
            10'd125: data <= 32'hfff5ff8d;
            10'd126: data <= 32'h001a0043;
            10'd127: data <= 32'h001a00ca;
            10'd128: data <= 32'hffb1005e;
            10'd129: data <= 32'hff75ffc7;
            10'd130: data <= 32'hff31ff2c;
            10'd131: data <= 32'hffde0062;
            10'd132: data <= 32'hff10ffbc;
            10'd133: data <= 32'hff5bffc1;
            10'd134: data <= 32'hff31ffcd;
            10'd135: data <= 32'hff580013;
            10'd136: data <= 32'hfeddff60;
            10'd137: data <= 32'hff88003f;
            10'd138: data <= 32'hff0f0000;
            10'd139: data <= 32'hfed1ff15;
            10'd140: data <= 32'hff810005;
            10'd141: data <= 32'hfee1ff60;
            10'd142: data <= 32'hff910003;
            10'd143: data <= 32'hff46fff3;
            10'd144: data <= 32'hff6affcd;
            10'd145: data <= 32'hff5bff91;
            10'd146: data <= 32'hfff3006c;
            10'd147: data <= 32'hff980018;
            10'd148: data <= 32'h002b00ab;
            10'd149: data <= 32'hff5aff58;
            10'd150: data <= 32'h003efff2;
            10'd151: data <= 32'hffe5ffc2;
            10'd152: data <= 32'h002bffb8;
            10'd153: data <= 32'h0026ffa1;
            10'd154: data <= 32'h00c80096;
            10'd155: data <= 32'h0036ffe5;
            10'd156: data <= 32'h00ed008b;
            10'd157: data <= 32'h008f004d;
            10'd158: data <= 32'h00e20072;
            10'd159: data <= 32'h00a10017;
            10'd160: data <= 32'h00b8ffe5;
            10'd161: data <= 32'h00a3ffac;
            10'd162: data <= 32'h00aeff97;
            10'd163: data <= 32'h007fff38;
            10'd164: data <= 32'h00d4ffad;
            10'd165: data <= 32'h0095ff94;
            10'd166: data <= 32'h00ceffe8;
            10'd167: data <= 32'h008fffcb;
            10'd168: data <= 32'h00a1ffe2;
            10'd169: data <= 32'h008cfffa;
            10'd170: data <= 32'h005fffca;
            10'd171: data <= 32'h0059ffce;
            10'd172: data <= 32'h0045ffe0;
            10'd173: data <= 32'h00a400d3;
            10'd174: data <= 32'hfff20032;
            10'd175: data <= 32'hffdcffa8;
            10'd176: data <= 32'h0021004c;
            10'd177: data <= 32'hff9bffd8;
            10'd178: data <= 32'hfff60052;
            10'd179: data <= 32'hff16ff37;
            10'd180: data <= 32'h005b0116;
            10'd181: data <= 32'hff6400ba;
            10'd182: data <= 32'hff46ffe7;
            10'd183: data <= 32'hff660015;
            10'd184: data <= 32'hff6b005d;
            10'd185: data <= 32'hfefbffaa;
            10'd186: data <= 32'hff7a0046;
            10'd187: data <= 32'hfef9ffce;
            10'd188: data <= 32'hffd90110;
            10'd189: data <= 32'hfeee0027;
            10'd190: data <= 32'hff33ffc2;
            10'd191: data <= 32'hff9a0096;
            10'd192: data <= 32'hff18ffe8;
            10'd193: data <= 32'hffdf00c8;
            10'd194: data <= 32'hff660073;
            10'd195: data <= 32'hff72ffe7;
            10'd196: data <= 32'h005d0172;
            10'd197: data <= 32'hff30ffdc;
            10'd198: data <= 32'h00020008;
            10'd199: data <= 32'hffaaffbc;
            10'd200: data <= 32'h0012ffe8;
            10'd201: data <= 32'h003b004d;
            10'd202: data <= 32'hff76feb1;
            10'd203: data <= 32'h00d10033;
            10'd204: data <= 32'h0008ffb6;
            10'd205: data <= 32'h00bf0031;
            10'd206: data <= 32'h005cffe2;
            10'd207: data <= 32'h00f60084;
            10'd208: data <= 32'h0078fff7;
            10'd209: data <= 32'h01550111;
            10'd210: data <= 32'h0049ffc3;
            10'd211: data <= 32'h00ff000a;
            10'd212: data <= 32'h00e40061;
            10'd213: data <= 32'h00afffee;
            10'd214: data <= 32'h00d50003;
            10'd215: data <= 32'h0090ffaa;
            10'd216: data <= 32'h00da0007;
            10'd217: data <= 32'h0075ffaa;
            10'd218: data <= 32'h0079ff7a;
            10'd219: data <= 32'h004bff45;
            10'd220: data <= 32'h0090ffd1;
            10'd221: data <= 32'h0061fffd;
            10'd222: data <= 32'hfff3ff47;
            10'd223: data <= 32'h0002ff31;
            10'd224: data <= 32'h004a0007;
            10'd225: data <= 32'hfffc0011;
            10'd226: data <= 32'hffe7fffd;
            10'd227: data <= 32'hffe4002c;
            10'd228: data <= 32'hffb20012;
            10'd229: data <= 32'hff6cff9e;
            10'd230: data <= 32'h000200bc;
            10'd231: data <= 32'hff630062;
            10'd232: data <= 32'hff24ff8e;
            10'd233: data <= 32'hff71fffa;
            10'd234: data <= 32'hff27ffd4;
            10'd235: data <= 32'hff2affb4;
            10'd236: data <= 32'hff33ffd9;
            10'd237: data <= 32'hff52002d;
            10'd238: data <= 32'hff280005;
            10'd239: data <= 32'hff02ff8e;
            10'd240: data <= 32'hff37ffb2;
            10'd241: data <= 32'hff9b008d;
            10'd242: data <= 32'hfebaff26;
            10'd243: data <= 32'hff32fefc;
            10'd244: data <= 32'hff2bff0c;
            10'd245: data <= 32'hff96ffa0;
            10'd246: data <= 32'hffa0ffed;
            10'd247: data <= 32'hfffc0083;
            10'd248: data <= 32'hffb4001a;
            10'd249: data <= 32'h000f0045;
            10'd250: data <= 32'hffe3fff6;
            10'd251: data <= 32'hffc6ff41;
            10'd252: data <= 32'h0029ff85;
            10'd253: data <= 32'h0038ffb4;
            10'd254: data <= 32'h004effb1;
            10'd255: data <= 32'h00af0049;
            10'd256: data <= 32'h005bffd4;
            10'd257: data <= 32'h00b0fff5;
            10'd258: data <= 32'h00b40019;
            10'd259: data <= 32'h00bb000d;
            10'd260: data <= 32'h00fa0074;
            10'd261: data <= 32'h007bffaa;
            10'd262: data <= 32'h00d2ffc1;
            10'd263: data <= 32'h00e20022;
            10'd264: data <= 32'h00eb0059;
            10'd265: data <= 32'h007effa6;
            10'd266: data <= 32'h00df0007;
            10'd267: data <= 32'h0063ff8a;
            10'd268: data <= 32'h00e00030;
            10'd269: data <= 32'h0046ffb0;
            10'd270: data <= 32'h004aff5d;
            10'd271: data <= 32'h008c000a;
            10'd272: data <= 32'h0036fff1;
            10'd273: data <= 32'h0026ffd0;
            10'd274: data <= 32'h000affce;
            10'd275: data <= 32'hfff8ffd6;
            10'd276: data <= 32'hffceffbb;
            10'd277: data <= 32'h003700af;
            10'd278: data <= 32'hff6bffe0;
            10'd279: data <= 32'hff54ff30;
            10'd280: data <= 32'hff75ff77;
            10'd281: data <= 32'hff7bffda;
            10'd282: data <= 32'hff98005f;
            10'd283: data <= 32'hff20ffd4;
            10'd284: data <= 32'hff33ffa9;
            10'd285: data <= 32'hff530007;
            10'd286: data <= 32'hff09ffb0;
            10'd287: data <= 32'hff500001;
            10'd288: data <= 32'hff1cffe5;
            10'd289: data <= 32'hff63003c;
            10'd290: data <= 32'hfee9ff84;
            10'd291: data <= 32'hff37ff85;
            10'd292: data <= 32'hff3effac;
            10'd293: data <= 32'hff940039;
            10'd294: data <= 32'hff64000d;
            10'd295: data <= 32'hff79ffd8;
            10'd296: data <= 32'hff8effcc;
            10'd297: data <= 32'hffcd0014;
            10'd298: data <= 32'hffd1001a;
            10'd299: data <= 32'h003600a9;
            10'd300: data <= 32'hfff10043;
            10'd301: data <= 32'h0063009c;
            10'd302: data <= 32'hffcdff94;
            10'd303: data <= 32'h005cffc2;
            10'd304: data <= 32'h0050ffde;
            10'd305: data <= 32'h009c002f;
            10'd306: data <= 32'h009f004c;
            10'd307: data <= 32'h0094000d;
            10'd308: data <= 32'h007fffa3;
            10'd309: data <= 32'h00a4ffa1;
            10'd310: data <= 32'h00c6ffe0;
            10'd311: data <= 32'h00f4004e;
            10'd312: data <= 32'h00ba000d;
            10'd313: data <= 32'h0094ff88;
            10'd314: data <= 32'h00f50015;
            10'd315: data <= 32'h00c10021;
            10'd316: data <= 32'h0066ff60;
            10'd317: data <= 32'h0085ff52;
            10'd318: data <= 32'h00d8002d;
            10'd319: data <= 32'h0093003b;
            10'd320: data <= 32'h00a30066;
            10'd321: data <= 32'h0011ff98;
            10'd322: data <= 32'h0026ff65;
            10'd323: data <= 32'h005f0019;
            10'd324: data <= 32'hffc6ff79;
            10'd325: data <= 32'h0023ffe7;
            10'd326: data <= 32'hffa0ff85;
            10'd327: data <= 32'hffc7ff9d;
            10'd328: data <= 32'hffabffcc;
            10'd329: data <= 32'hff6eff86;
            10'd330: data <= 32'hffc30031;
            10'd331: data <= 32'hff3dffc4;
            10'd332: data <= 32'hff61ffc2;
            10'd333: data <= 32'hff13ff6e;
            10'd334: data <= 32'hffce00b7;
            10'd335: data <= 32'hff4c00a5;
            10'd336: data <= 32'hfef1ffa6;
            10'd337: data <= 32'hff41ffda;
            10'd338: data <= 32'hff770087;
            10'd339: data <= 32'hff6200a1;
            10'd340: data <= 32'hff1a0002;
            10'd341: data <= 32'hff3affd5;
            10'd342: data <= 32'hff2aff9d;
            10'd343: data <= 32'hffcc009c;
            10'd344: data <= 32'hff4d0021;
            10'd345: data <= 32'hff9a0011;
            10'd346: data <= 32'hffaf0039;
            10'd347: data <= 32'hffc8003e;
            10'd348: data <= 32'hff8aff98;
            10'd349: data <= 32'h0000ffee;
            10'd350: data <= 32'hfffe0009;
            10'd351: data <= 32'hffd8ff79;
            10'd352: data <= 32'h0009ff5d;
            10'd353: data <= 32'h005effdf;
            10'd354: data <= 32'h00850044;
            10'd355: data <= 32'h00bf00b3;
            10'd356: data <= 32'h0038ffb8;
            10'd357: data <= 32'h0099ffae;
            10'd358: data <= 32'h00d6003e;
            10'd359: data <= 32'h00b80027;
            10'd360: data <= 32'h00b2ffe9;
            10'd361: data <= 32'h0105006c;
            10'd362: data <= 32'h00a8fffe;
            10'd363: data <= 32'h00a3ff95;
            10'd364: data <= 32'h00c3ffc1;
            10'd365: data <= 32'h00b6ffd1;
            10'd366: data <= 32'h01000075;
            10'd367: data <= 32'hffebfec9;
            10'd368: data <= 32'h00f5ffd8;
            10'd369: data <= 32'h00ce00b8;
            10'd370: data <= 32'h0042ffe7;
            10'd371: data <= 32'h0061ffd4;
            10'd372: data <= 32'h00b000c2;
            10'd373: data <= 32'hfff1ffef;
            10'd374: data <= 32'hfffcff93;
            10'd375: data <= 32'hffd4ff7e;
            10'd376: data <= 32'hfffcffe7;
            10'd377: data <= 32'hffa6ffb5;
            10'd378: data <= 32'hff77ff53;
            10'd379: data <= 32'hff80ff6c;
            10'd380: data <= 32'hffed008a;
            10'd381: data <= 32'hff3bfff0;
            10'd382: data <= 32'hffb50075;
            10'd383: data <= 32'hfeedff8e;
            10'd384: data <= 32'hff5effc8;
            10'd385: data <= 32'hff3b0000;
            10'd386: data <= 32'hff2dffe7;
            10'd387: data <= 32'hfef1ff6d;
            10'd388: data <= 32'hff4dffde;
            10'd389: data <= 32'hff9900c9;
            10'd390: data <= 32'hfeb6ff63;
            10'd391: data <= 32'hffa40035;
            10'd392: data <= 32'hff16ffd8;
            10'd393: data <= 32'hff03ff05;
            10'd394: data <= 32'hffda004b;
            10'd395: data <= 32'hff7b003c;
            10'd396: data <= 32'hff93ffea;
            10'd397: data <= 32'hff86ff99;
            10'd398: data <= 32'h00030031;
            10'd399: data <= 32'hffbcffd9;
            10'd400: data <= 32'hfffcffce;
            10'd401: data <= 32'h004a0053;
            10'd402: data <= 32'h001a0002;
            10'd403: data <= 32'h004affed;
            10'd404: data <= 32'h005efff6;
            10'd405: data <= 32'h00d000aa;
            10'd406: data <= 32'h00720035;
            10'd407: data <= 32'h00a4000b;
            10'd408: data <= 32'h00ca0049;
            10'd409: data <= 32'h00e60081;
            10'd410: data <= 32'h00aa0011;
            10'd411: data <= 32'h01070075;
            10'd412: data <= 32'h00d5005e;
            10'd413: data <= 32'h0093ffad;
            10'd414: data <= 32'h017d0131;
            10'd415: data <= 32'h0014ff71;
            10'd416: data <= 32'h0115001b;
            10'd417: data <= 32'h006cffd0;
            10'd418: data <= 32'h009effc2;
            10'd419: data <= 32'h006cffb4;
            10'd420: data <= 32'h008d0000;
            10'd421: data <= 32'h003bffbd;
            10'd422: data <= 32'h004fffd9;
            10'd423: data <= 32'h0030fff3;
            10'd424: data <= 32'h0024000c;
            10'd425: data <= 32'hffd9ffba;
            10'd426: data <= 32'h001f0045;
            10'd427: data <= 32'hffa5ffe8;
            10'd428: data <= 32'hff58ff23;
            10'd429: data <= 32'hffe40015;
            10'd430: data <= 32'hffa5006d;
            10'd431: data <= 32'hff7c0038;
            10'd432: data <= 32'hff4bffe8;
            10'd433: data <= 32'hffab009b;
            10'd434: data <= 32'hfed1ff78;
            10'd435: data <= 32'hff46ff9e;
            10'd436: data <= 32'hff3cfffc;
            10'd437: data <= 32'hff520039;
            10'd438: data <= 32'hff70009a;
            10'd439: data <= 32'hfec2ff68;
            10'd440: data <= 32'hffbb0084;
            10'd441: data <= 32'hff240035;
            10'd442: data <= 32'hff57fff8;
            10'd443: data <= 32'hff31ffa3;
            10'd444: data <= 32'hff7bffd5;
            10'd445: data <= 32'hff47ff77;
            10'd446: data <= 32'hffdf002f;
            10'd447: data <= 32'hff7fffcb;
            10'd448: data <= 32'hffcaffc2;
            10'd449: data <= 32'hffc0ffa1;
            10'd450: data <= 32'hfffaffbd;
            10'd451: data <= 32'h0014ffde;
            10'd452: data <= 32'hfff2ff6e;
            10'd453: data <= 32'h0084001c;
            10'd454: data <= 32'h00680038;
            10'd455: data <= 32'h00bc0095;
            10'd456: data <= 32'h00be00bb;
            10'd457: data <= 32'h007b000f;
            10'd458: data <= 32'h00d3003e;
            10'd459: data <= 32'h004eff5a;
            10'd460: data <= 32'h00cbff9f;
            10'd461: data <= 32'h00c3ffe5;
            10'd462: data <= 32'h008fff77;
            10'd463: data <= 32'h00c5ffa3;
            10'd464: data <= 32'h00ee002c;
            10'd465: data <= 32'h00bc0011;
            10'd466: data <= 32'h012a00de;
            10'd467: data <= 32'h00830034;
            10'd468: data <= 32'h00c3003b;
            10'd469: data <= 32'h007a000c;
            10'd470: data <= 32'h0039ff7a;
            10'd471: data <= 32'h0074ffda;
            10'd472: data <= 32'h008d0088;
            10'd473: data <= 32'hffc0ff66;
            10'd474: data <= 32'h006f0034;
            10'd475: data <= 32'hfff40030;
            10'd476: data <= 32'hff80ff30;
            10'd477: data <= 32'h00410070;
            10'd478: data <= 32'hffc30089;
            10'd479: data <= 32'hffc70078;
            10'd480: data <= 32'hff21ff74;
            10'd481: data <= 32'hffbe002c;
            10'd482: data <= 32'hff63003f;
            10'd483: data <= 32'hff93008d;
            10'd484: data <= 32'hff0affdb;
            10'd485: data <= 32'hffa10095;
            10'd486: data <= 32'hff050009;
            10'd487: data <= 32'hfed0ff18;
            10'd488: data <= 32'hff8c0036;
            10'd489: data <= 32'hfef6ffc7;
            10'd490: data <= 32'hff5f0001;
            10'd491: data <= 32'hff640054;
            10'd492: data <= 32'hff90009e;
            10'd493: data <= 32'hff2fffeb;
            10'd494: data <= 32'hff1dff2c;
            10'd495: data <= 32'hffb4ffe9;
            10'd496: data <= 32'hff9a000d;
            10'd497: data <= 32'hff90ffb2;
            10'd498: data <= 32'hffe30000;
            10'd499: data <= 32'h003700b0;
            10'd500: data <= 32'hffc8fff0;
            10'd501: data <= 32'hfff7ff90;
            10'd502: data <= 32'h008b0080;
            10'd503: data <= 32'h0002ffc9;
            10'd504: data <= 32'h00bb006f;
            10'd505: data <= 32'h0060002f;
            10'd506: data <= 32'h00a4002a;
            10'd507: data <= 32'h008cffff;
            10'd508: data <= 32'h00a3ffe4;
            10'd509: data <= 32'h00afffe1;
            10'd510: data <= 32'h0099ff9f;
            10'd511: data <= 32'h00b1ff9b;
            10'd512: data <= 32'h00e40005;
            10'd513: data <= 32'h00cd0010;
            10'd514: data <= 32'h00a6ffbe;
            10'd515: data <= 32'h008bff69;
            10'd516: data <= 32'h00c6ffcd;
            10'd517: data <= 32'h009dffda;
            10'd518: data <= 32'h0046ff3a;
            10'd519: data <= 32'h009effb5;
            10'd520: data <= 32'h0073ffed;
            10'd521: data <= 32'h0070000b;
            10'd522: data <= 32'h008b008a;
            10'd523: data <= 32'hffebffbd;
            10'd524: data <= 32'h000bffa0;
            10'd525: data <= 32'h0025002b;
            10'd526: data <= 32'hffafffb3;
            10'd527: data <= 32'hfff2000e;
            10'd528: data <= 32'hffb20019;
            10'd529: data <= 32'hff41ff47;
            10'd530: data <= 32'h00020086;
            10'd531: data <= 32'hff420010;
            10'd532: data <= 32'hff43ff9e;
            10'd533: data <= 32'hffb900a0;
            10'd534: data <= 32'hff420061;
            10'd535: data <= 32'hff42001b;
            10'd536: data <= 32'hff23ffe9;
            10'd537: data <= 32'hff26ffd1;
            10'd538: data <= 32'hff2cffda;
            10'd539: data <= 32'hff9500ad;
            10'd540: data <= 32'hfefaffe5;
            10'd541: data <= 32'hff68000b;
            10'd542: data <= 32'hff72005a;
            10'd543: data <= 32'hff0dff7f;
            10'd544: data <= 32'hff6fff9c;
            10'd545: data <= 32'hfff100b7;
            10'd546: data <= 32'hff9f0074;
            10'd547: data <= 32'hffe3007a;
            10'd548: data <= 32'hff9effe7;
            10'd549: data <= 32'h00130034;
            10'd550: data <= 32'hffcfffcd;
            10'd551: data <= 32'h004b0035;
            10'd552: data <= 32'h0004ffd6;
            10'd553: data <= 32'h0088004e;
            10'd554: data <= 32'h0069004d;
            10'd555: data <= 32'h0057ffd6;
            10'd556: data <= 32'h010d00e4;
            10'd557: data <= 32'h0062001e;
            10'd558: data <= 32'h006eff62;
            10'd559: data <= 32'h00cbffd9;
            10'd560: data <= 32'h005bff34;
            10'd561: data <= 32'h012d0048;
            10'd562: data <= 32'h008effdc;
            10'd563: data <= 32'h011f006b;
            10'd564: data <= 32'h0078ffb6;
            10'd565: data <= 32'h00fe0029;
            10'd566: data <= 32'h0094ffed;
            10'd567: data <= 32'h0088ff97;
            10'd568: data <= 32'h00b70001;
            10'd569: data <= 32'h00aa004e;
            10'd570: data <= 32'h0059ffe9;
            10'd571: data <= 32'h007a0016;
            10'd572: data <= 32'h0000ff7f;
            10'd573: data <= 32'h002aff99;
            10'd574: data <= 32'h0009ffc1;
            10'd575: data <= 32'hfffbffd6;
            10'd576: data <= 32'h002f0080;
            10'd577: data <= 32'hffbf0033;
            10'd578: data <= 32'hffb0fff8;
            10'd579: data <= 32'hffdf007f;
            10'd580: data <= 32'hff81003f;
            10'd581: data <= 32'hff47ffb2;
            10'd582: data <= 32'hffb50076;
            10'd583: data <= 32'hff330016;
            10'd584: data <= 32'hff3effdc;
            10'd585: data <= 32'hff650044;
            10'd586: data <= 32'hff230004;
            10'd587: data <= 32'hff650054;
            10'd588: data <= 32'hff590085;
            10'd589: data <= 32'hfee1ff90;
            10'd590: data <= 32'hfeecff08;
            10'd591: data <= 32'hff7ffffb;
            10'd592: data <= 32'hff3efff5;
            10'd593: data <= 32'hff9a0056;
            10'd594: data <= 32'hff680025;
            10'd595: data <= 32'hff27ff3d;
            10'd596: data <= 32'hfff10032;
            10'd597: data <= 32'hff53ff82;
            10'd598: data <= 32'hffc9ff8f;
            10'd599: data <= 32'hfff80004;
            10'd600: data <= 32'hffc5ff91;
            10'd601: data <= 32'hffbafef6;
            10'd602: data <= 32'h009b004a;
            10'd603: data <= 32'hffbeff38;
            10'd604: data <= 32'h00affffc;
            10'd605: data <= 32'h0074002d;
            10'd606: data <= 32'h0082ffee;
            10'd607: data <= 32'h00b9002c;
            10'd608: data <= 32'h00ba0039;
            10'd609: data <= 32'h008effc0;
            10'd610: data <= 32'h010f006d;
            10'd611: data <= 32'h0094ffe8;
            10'd612: data <= 32'h00ff0039;
            10'd613: data <= 32'h00c90030;
            10'd614: data <= 32'h00eb004e;
            10'd615: data <= 32'h00f60094;
            10'd616: data <= 32'h007effd6;
            10'd617: data <= 32'h00a8ffc7;
            10'd618: data <= 32'h00b70026;
            10'd619: data <= 32'h007e0000;
            10'd620: data <= 32'h00bf0085;
            10'd621: data <= 32'h0032fff5;
            10'd622: data <= 32'h0000ff46;
            10'd623: data <= 32'h0047ffca;
            10'd624: data <= 32'hffb0ff2b;
            10'd625: data <= 32'h00430002;
            10'd626: data <= 32'hffbbffd7;
            10'd627: data <= 32'hffbeffb0;
            10'd628: data <= 32'hffc80005;
            10'd629: data <= 32'hff4eff6d;
            10'd630: data <= 32'hffe10051;
            10'd631: data <= 32'hff670036;
            10'd632: data <= 32'hff39ffad;
            10'd633: data <= 32'hff4affbe;
            10'd634: data <= 32'hff4dfff5;
            10'd635: data <= 32'hff720065;
            10'd636: data <= 32'hfea9ff20;
            10'd637: data <= 32'hff80fffe;
            10'd638: data <= 32'hfee3ff93;
            10'd639: data <= 32'hff6a0009;
            10'd640: data <= 32'hff50004a;
            10'd641: data <= 32'hfebaff02;
            10'd642: data <= 32'hffac000e;
            10'd643: data <= 32'hff42ffff;
            10'd644: data <= 32'hff74ffe1;
            10'd645: data <= 32'hff6bffc0;
            10'd646: data <= 32'hffb8000d;
            10'd647: data <= 32'hff61ff69;
            10'd648: data <= 32'hffbfff81;
            10'd649: data <= 32'hffa6ff54;
            10'd650: data <= 32'h002afff6;
            10'd651: data <= 32'hffefffc1;
            10'd652: data <= 32'h0007ff76;
            10'd653: data <= 32'h0083002d;
            10'd654: data <= 32'h007e0066;
            10'd655: data <= 32'h00750022;
            10'd656: data <= 32'h007bffe9;
            10'd657: data <= 32'h00ae0012;
            10'd658: data <= 32'h008dffd2;
            10'd659: data <= 32'h00b5ffd8;
            10'd660: data <= 32'h0096ff9d;
            10'd661: data <= 32'h00e4fffe;
            10'd662: data <= 32'h012e00d5;
            10'd663: data <= 32'h00e0009e;
            10'd664: data <= 32'h00be0021;
            10'd665: data <= 32'h01070091;
            10'd666: data <= 32'h00bc005d;
            10'd667: data <= 32'h008fffe3;
            10'd668: data <= 32'h00db0067;
            10'd669: data <= 32'h006d000a;
            10'd670: data <= 32'h00a8004d;
            10'd671: data <= 32'h007d006e;
            10'd672: data <= 32'h0049002b;
            10'd673: data <= 32'hfff8ff98;
            10'd674: data <= 32'h007f008d;
            10'd675: data <= 32'hff9effa6;
            10'd676: data <= 32'h001b000c;
            10'd677: data <= 32'hffb3fff9;
            10'd678: data <= 32'hff8cff97;
            10'd679: data <= 32'hff8affa3;
            10'd680: data <= 32'hffa1000b;
            10'd681: data <= 32'hff2cff80;
            10'd682: data <= 32'hff82ffea;
            10'd683: data <= 32'hff3bffde;
            10'd684: data <= 32'hff50fff3;
            10'd685: data <= 32'hff660053;
            10'd686: data <= 32'hff11ffe2;
            10'd687: data <= 32'hff5e0031;
            10'd688: data <= 32'hff10ffe3;
            10'd689: data <= 32'hff48ffff;
            10'd690: data <= 32'hff03ff97;
            10'd691: data <= 32'hff840034;
            10'd692: data <= 32'hff36fffc;
            10'd693: data <= 32'hff6bfff8;
            10'd694: data <= 32'hffde00d9;
            10'd695: data <= 32'hff23ffb5;
            10'd696: data <= 32'hffce0006;
            10'd697: data <= 32'hff84ffc7;
            10'd698: data <= 32'h005200d7;
            10'd699: data <= 32'hff88ffd7;
            10'd700: data <= 32'h0043003b;
            10'd701: data <= 32'hffdbffc5;
            10'd702: data <= 32'h0034ffc6;
            10'd703: data <= 32'h0027ffae;
            10'd704: data <= 32'h0034ff75;
            10'd705: data <= 32'h00ab0020;
            10'd706: data <= 32'h0052ffb6;
            10'd707: data <= 32'h009dffc0;
            10'd708: data <= 32'h00f70084;
            10'd709: data <= 32'h00ac0036;
            10'd710: data <= 32'h00f6006a;
            10'd711: data <= 32'h0066ff7f;
            10'd712: data <= 32'h0104000c;
            10'd713: data <= 32'h00c00015;
            10'd714: data <= 32'h009dffa3;
            10'd715: data <= 32'h00c4ffcf;
            10'd716: data <= 32'h00bcfffb;
            10'd717: data <= 32'h00b00003;
            10'd718: data <= 32'h00aa001c;
            10'd719: data <= 32'h0030ff58;
            10'd720: data <= 32'h006cff7d;
            10'd721: data <= 32'hfffeff0b;
            10'd722: data <= 32'h00c10060;
            10'd723: data <= 32'hffc8ff8f;
            10'd724: data <= 32'h003effdd;
            10'd725: data <= 32'hffa5ff5c;
            10'd726: data <= 32'h0004ffcc;
            10'd727: data <= 32'hffb5ffd4;
            10'd728: data <= 32'hffbbffea;
            10'd729: data <= 32'hff41ff43;
            10'd730: data <= 32'h001100a0;
            10'd731: data <= 32'hff02ffa0;
            10'd732: data <= 32'hff76ffba;
            10'd733: data <= 32'hff0bff6f;
            10'd734: data <= 32'hff40ff94;
            10'd735: data <= 32'hff980091;
            10'd736: data <= 32'hfef1ffd2;
            10'd737: data <= 32'hff6e0034;
            10'd738: data <= 32'hff5f008e;
            10'd739: data <= 32'hff250019;
            10'd740: data <= 32'hff0bff97;
            10'd741: data <= 32'hff9a006b;
            10'd742: data <= 32'hff23fff2;
            10'd743: data <= 32'hffa20057;
            10'd744: data <= 32'hff2effbb;
            10'd745: data <= 32'hffdc0064;
            10'd746: data <= 32'hffad0073;
            10'd747: data <= 32'hff7cffb5;
            10'd748: data <= 32'hffc2ffb4;
            10'd749: data <= 32'hff97ff48;
            10'd750: data <= 32'h004d0031;
            10'd751: data <= 32'hffefffea;
            10'd752: data <= 32'h002fffd2;
            10'd753: data <= 32'h00ad00b8;
            10'd754: data <= 32'h001dffe6;
            10'd755: data <= 32'h011e0114;
            10'd756: data <= 32'h00470034;
            10'd757: data <= 32'h00c00022;
            10'd758: data <= 32'h00d6007d;
            10'd759: data <= 32'h0071ffaf;
            10'd760: data <= 32'h00c3ffbe;
            10'd761: data <= 32'h00e70030;
            10'd762: data <= 32'h0099ffb9;
            10'd763: data <= 32'h0106003e;
            10'd764: data <= 32'h0096ffd4;
            10'd765: data <= 32'h00f00029;
            10'd766: data <= 32'h00f1009b;
            10'd767: data <= 32'h00920018;
            10'd768: data <= 32'h009efff8;
            10'd769: data <= 32'h00e000ab;
            10'd770: data <= 32'h004a0009;
            10'd771: data <= 32'h00730005;
            10'd772: data <= 32'h003dfff9;
            10'd773: data <= 32'h0038ffff;
            10'd774: data <= 32'h0007ffe0;
            10'd775: data <= 32'hffb3ff52;
            10'd776: data <= 32'hffcfff6e;
            10'd777: data <= 32'h00190060;
            10'd778: data <= 32'hff80ffdd;
            10'd779: data <= 32'hfffd008e;
            10'd780: data <= 32'hffd000f7;
            10'd781: data <= 32'hff84008d;
            10'd782: data <= 32'hfef3ff56;
            10'd783: data <= 32'hffbe0064;
            10'd784: data <= 32'hfeaeff32;
            10'd785: data <= 32'hff70ffc4;
            10'd786: data <= 32'hff4e0045;
            10'd787: data <= 32'hff530057;
            10'd788: data <= 32'hfec8ff53;
            10'd789: data <= 32'hff70fffd;
            10'd790: data <= 32'hff9300d0;
            10'd791: data <= 32'hfee2ffa1;
            10'd792: data <= 32'hff55ffa9;
            10'd793: data <= 32'hff40ffab;
            10'd794: data <= 32'hffcd007e;
            10'd795: data <= 32'hff49ffde;
            10'd796: data <= 32'hff7dff89;
            10'd797: data <= 32'hffeb0038;
            10'd798: data <= 32'hffc5001e;
            10'd799: data <= 32'hffdbffe9;
            10'd800: data <= 32'hffb8ff65;
            10'd801: data <= 32'h0040fff4;
            10'd802: data <= 32'h001cffea;
            10'd803: data <= 32'h00a7009e;
            10'd804: data <= 32'h005e0060;
            10'd805: data <= 32'h00c800b5;
            10'd806: data <= 32'h0046ffdf;
            10'd807: data <= 32'h00c30014;
            10'd808: data <= 32'h00f000ab;
            10'd809: data <= 32'h007cffe1;
            10'd810: data <= 32'h009eff89;
            10'd811: data <= 32'h00defffa;
            10'd812: data <= 32'h007cff6b;
            10'd813: data <= 32'h00ceffa5;
            10'd814: data <= 32'h008eff77;
            10'd815: data <= 32'h00ff0027;
            10'd816: data <= 32'h00a30004;
            10'd817: data <= 32'h005aff4a;
            10'd818: data <= 32'h013300c4;
            10'd819: data <= 32'h0005ff89;
            10'd820: data <= 32'h0093ffb6;
            10'd821: data <= 32'h00790034;
            10'd822: data <= 32'h0015ffac;
            10'd823: data <= 32'h0000ff5d;
            10'd824: data <= 32'hfff3ff67;
            10'd825: data <= 32'h00450043;
            10'd826: data <= 32'h000d0089;
            10'd827: data <= 32'hffd6004b;
            10'd828: data <= 32'hff6dff8c;
            10'd829: data <= 32'hffcd0011;
            10'd830: data <= 32'hff970043;
            10'd831: data <= 32'hff680001;
            10'd832: data <= 32'hff6d0010;
            10'd833: data <= 32'hff48fff7;
            10'd834: data <= 32'hff55000f;
            10'd835: data <= 32'hff31fff5;
            10'd836: data <= 32'hff7a0079;
            10'd837: data <= 32'hfecfff84;
            10'd838: data <= 32'hff8a0046;
            10'd839: data <= 32'hff380051;
            10'd840: data <= 32'hff31fff8;
            10'd841: data <= 32'hff43fff2;
            10'd842: data <= 32'hff50fff5;
            10'd843: data <= 32'hff720018;
            10'd844: data <= 32'hffa80079;
            10'd845: data <= 32'hff64fffb;
            10'd846: data <= 32'hff79ff9f;
            10'd847: data <= 32'hff97ff95;
            10'd848: data <= 32'hfffb0029;
            10'd849: data <= 32'h0008006a;
            10'd850: data <= 32'hffe6fffc;
            10'd851: data <= 32'h00340024;
            10'd852: data <= 32'h007700a6;
            10'd853: data <= 32'h00320026;
            10'd854: data <= 32'h005efff3;
            10'd855: data <= 32'h0039ff82;
            10'd856: data <= 32'h0080ff9e;
            10'd857: data <= 32'h00e00063;
            10'd858: data <= 32'h0082ffef;
            10'd859: data <= 32'h008cff84;
            10'd860: data <= 32'h01220082;
            10'd861: data <= 32'h007affc4;
            10'd862: data <= 32'h00eefffc;
            10'd863: data <= 32'h00c30009;
            10'd864: data <= 32'h00a6ffb3;
            10'd865: data <= 32'h01140077;
            10'd866: data <= 32'h00cc007d;
            10'd867: data <= 32'h0048ff63;
            10'd868: data <= 32'h0051feff;
            10'd869: data <= 32'h01030078;
            10'd870: data <= 32'h00830080;
            10'd871: data <= 32'h005e001b;
            10'd872: data <= 32'hfffaff67;
            10'd873: data <= 32'h007c0035;
            10'd874: data <= 32'h0000000a;
            10'd875: data <= 32'h001f002d;
            10'd876: data <= 32'h00000057;
            10'd877: data <= 32'hff5cff45;
            10'd878: data <= 32'hffc7ffa8;
            10'd879: data <= 32'h000000bd;
            10'd880: data <= 32'hff830064;
            10'd881: data <= 32'hfee7fefd;
            10'd882: data <= 32'hff92ffc3;
            10'd883: data <= 32'hff500007;
            10'd884: data <= 32'hff44fff1;
            10'd885: data <= 32'hff780070;
            10'd886: data <= 32'hff7700c2;
            10'd887: data <= 32'hfedeffaf;
            10'd888: data <= 32'hff8b0062;
            10'd889: data <= 32'hfed0ff8c;
            10'd890: data <= 32'hffae0079;
            10'd891: data <= 32'hff180013;
            10'd892: data <= 32'hff20ff7b;
            10'd893: data <= 32'hff6effd6;
            10'd894: data <= 32'hff9e004f;
            10'd895: data <= 32'hff6ffffb;
            10'd896: data <= 32'hff9cffeb;
            10'd897: data <= 32'hffa6ffdd;
            10'd898: data <= 32'hffb0ffb1;
            10'd899: data <= 32'h0000000c;
            10'd900: data <= 32'h00270063;
            10'd901: data <= 32'h0027004c;
            10'd902: data <= 32'h000bffcf;
            10'd903: data <= 32'h0074002d;
            10'd904: data <= 32'h001cff9e;
            10'd905: data <= 32'h0087ffd4;
            10'd906: data <= 32'h005fffa7;
            10'd907: data <= 32'h012e00e7;
            10'd908: data <= 32'h0036ffb1;
            10'd909: data <= 32'h00f2000a;
            10'd910: data <= 32'h00ea007e;
            10'd911: data <= 32'h00a2ffeb;
            10'd912: data <= 32'h00e70018;
            10'd913: data <= 32'h00f80074;
            10'd914: data <= 32'h00d70056;
            10'd915: data <= 32'h00b40006;
            10'd916: data <= 32'h0081ff8f;
            10'd917: data <= 32'h009fffa4;
            10'd918: data <= 32'h00d30049;
            10'd919: data <= 32'h008d0037;
            10'd920: data <= 32'h0079000f;
            10'd921: data <= 32'h00680011;
            10'd922: data <= 32'h002affc7;
            10'd923: data <= 32'h002affcb;
            10'd924: data <= 32'h00340022;
            10'd925: data <= 32'h00050025;
            10'd926: data <= 32'hfffe003b;
            10'd927: data <= 32'hff90ffa6;
            10'd928: data <= 32'hff9eff92;
            10'd929: data <= 32'hff58ff49;
            10'd930: data <= 32'hff82ff91;
            10'd931: data <= 32'hff74ffdc;
            10'd932: data <= 32'hff89003c;
            10'd933: data <= 32'hff23ffc4;
            10'd934: data <= 32'hff87004c;
            10'd935: data <= 32'hff0fffe3;
            10'd936: data <= 32'hff3dffe1;
            10'd937: data <= 32'hff680065;
            10'd938: data <= 32'hff7700c1;
            10'd939: data <= 32'hfeefffcf;
            10'd940: data <= 32'hff4cffe4;
            10'd941: data <= 32'hff58002a;
            10'd942: data <= 32'hff88007c;
            10'd943: data <= 32'hff26ffcd;
            10'd944: data <= 32'hffa70031;
            10'd945: data <= 32'hffbe009f;
            10'd946: data <= 32'hff86001d;
            10'd947: data <= 32'hff9cffca;
            10'd948: data <= 32'hfff0002b;
            10'd949: data <= 32'hffa9ffa7;
            10'd950: data <= 32'h001afff3;
            10'd951: data <= 32'hffedffb7;
            10'd952: data <= 32'h0030ffc6;
            10'd953: data <= 32'h00860063;
            10'd954: data <= 32'h0035ffe5;
            10'd955: data <= 32'h0022ff2c;
            10'd956: data <= 32'h0099ffad;
            10'd957: data <= 32'h00c5003f;
            10'd958: data <= 32'h00b2002f;
            10'd959: data <= 32'h00da0051;
            10'd960: data <= 32'h00f70096;
            10'd961: data <= 32'h0143013f;
            10'd962: data <= 32'h00a10052;
            10'd963: data <= 32'h01050070;
            10'd964: data <= 32'h00cd0056;
            10'd965: data <= 32'h00b2fffb;
            10'd966: data <= 32'h008bff9f;
            10'd967: data <= 32'h00e90046;
            10'd968: data <= 32'h009a0035;
            10'd969: data <= 32'h00980023;
            10'd970: data <= 32'h0058ffd5;
            10'd971: data <= 32'h005dffd6;
            10'd972: data <= 32'h0003ff64;
            10'd973: data <= 32'h001cff7a;
            10'd974: data <= 32'h00460025;
            10'd975: data <= 32'h00080033;
            10'd976: data <= 32'h0023008a;
            10'd977: data <= 32'hffbf0032;
            10'd978: data <= 32'hff2ffef8;
            10'd979: data <= 32'hff89ff3b;
            10'd980: data <= 32'hff9fffec;
            10'd981: data <= 32'hff6dfff3;
            10'd982: data <= 32'hff52ffd2;
            10'd983: data <= 32'hff19ff73;
            10'd984: data <= 32'hff9e005e;
            10'd985: data <= 32'hfef0ffb5;
            10'd986: data <= 32'hff9e007f;
            10'd987: data <= 32'hff110024;
            10'd988: data <= 32'hff37fff5;
            10'd989: data <= 32'hff33fffb;
            10'd990: data <= 32'hff620044;
            10'd991: data <= 32'hff4b0031;
            10'd992: data <= 32'hffa100ab;
            10'd993: data <= 32'hff25ffe9;
            10'd994: data <= 32'hff5bffa0;
            10'd995: data <= 32'hff7affbf;
            10'd996: data <= 32'hffc1002b;
            10'd997: data <= 32'hff82ffbd;
            10'd998: data <= 32'hff88ff40;
            10'd999: data <= 32'h007900c6;
            10'd1000: data <= 32'hffc90024;
            10'd1001: data <= 32'h00660079;
            10'd1002: data <= 32'hffe3ffbc;
            10'd1003: data <= 32'h0045ffab;
            10'd1004: data <= 32'h005effe1;
            10'd1005: data <= 32'h00880013;
            10'd1006: data <= 32'h007bffed;
            10'd1007: data <= 32'h006cff8d;
            10'd1008: data <= 32'h00aaffbb;
            10'd1009: data <= 32'h00b8ffe8;
            10'd1010: data <= 32'h00c6fffd;
            10'd1011: data <= 32'h0075ff58;
            10'd1012: data <= 32'h00f3ffe8;
            10'd1013: data <= 32'h009affaf;
            10'd1014: data <= 32'h011a0065;
            10'd1015: data <= 32'h00ad0026;
            10'd1016: data <= 32'h00acffe0;
            10'd1017: data <= 32'h0071ff7b;
            10'd1018: data <= 32'h0099ffac;
            10'd1019: data <= 32'h00f800be;
            10'd1020: data <= 32'hfff6ff73;
            10'd1021: data <= 32'h00e50086;
            10'd1022: data <= 32'h00330051;
            10'd1023: data <= 32'h0049002a;
            default: data <= 32'h00000000;
        endcase
    end
endmodule
